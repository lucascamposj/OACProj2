library verilog;
use verilog.vl_types.all;
entity controlPC_vlg_vec_tst is
end controlPC_vlg_vec_tst;

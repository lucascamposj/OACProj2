library verilog;
use verilog.vl_types.all;
entity lui32_vlg_vec_tst is
end lui32_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity PipelineInit_vlg_vec_tst is
end PipelineInit_vlg_vec_tst;

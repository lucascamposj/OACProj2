library verilog;
use verilog.vl_types.all;
entity ShiftLeft_vlg_vec_tst is
end ShiftLeft_vlg_vec_tst;

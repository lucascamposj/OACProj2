library verilog;
use verilog.vl_types.all;
entity Equal5_vlg_vec_tst is
end Equal5_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity EXMEM_vlg_vec_tst is
end EXMEM_vlg_vec_tst;

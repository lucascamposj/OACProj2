library verilog;
use verilog.vl_types.all;
entity mux4to2_vlg_vec_tst is
end mux4to2_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity ShiftLeft2_vlg_vec_tst is
end ShiftLeft2_vlg_vec_tst;

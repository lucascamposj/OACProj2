library verilog;
use verilog.vl_types.all;
entity plusFour32_vlg_vec_tst is
end plusFour32_vlg_vec_tst;

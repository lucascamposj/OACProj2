library verilog;
use verilog.vl_types.all;
entity SignExtent_vlg_vec_tst is
end SignExtent_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity PipelineInit_vlg_check_tst is
    port(
        ALUOperation    : in     vl_logic_vector(3 downto 0);
        BInstruction    : in     vl_logic_vector(31 downto 0);
        BPC             : in     vl_logic_vector(31 downto 0);
        BproxPC         : in     vl_logic_vector(31 downto 0);
        DCtrlBranch     : in     vl_logic_vector(1 downto 0);
        DCtrlcontrolJump: in     vl_logic_vector(1 downto 0);
        DCtrlEscreveMem : in     vl_logic;
        DCtrlEscreveReg : in     vl_logic;
        DCtrlExtent     : in     vl_logic;
        DCtrlMemParaReg : in     vl_logic;
        DCtrlopALU      : in     vl_logic_vector(2 downto 0);
        DCtrlOrigALU    : in     vl_logic;
        DCtrlRegDst     : in     vl_logic_vector(1 downto 0);
        DInstruction    : in     vl_logic_vector(31 downto 0);
        DJAL            : in     vl_logic;
        DJump           : in     vl_logic;
        DJumpPC         : in     vl_logic_vector(31 downto 0);
        DRSDados0       : in     vl_logic_vector(31 downto 0);
        DRTDados1       : in     vl_logic_vector(31 downto 0);
        EXBranch        : in     vl_logic_vector(1 downto 0);
        EXHIGH          : in     vl_logic_vector(31 downto 0);
        EXImm           : in     vl_logic_vector(5 downto 0);
        EXLOW           : in     vl_logic_vector(31 downto 0);
        EXopALU         : in     vl_logic_vector(2 downto 0);
        EXULAA          : in     vl_logic_vector(31 downto 0);
        EXULAB          : in     vl_logic_vector(31 downto 0);
        Flush           : in     vl_logic;
        ForwardA        : in     vl_logic_vector(1 downto 0);
        ForwardB        : in     vl_logic_vector(1 downto 0);
        Jump            : in     vl_logic;
        MEMBranch       : in     vl_logic_vector(1 downto 0);
        MEMEscreveMem   : in     vl_logic;
        MEMnPC          : in     vl_logic_vector(31 downto 0);
        MEMReadValue    : in     vl_logic_vector(31 downto 0);
        MEMZero         : in     vl_logic;
        OrigPC          : in     vl_logic;
        outALU          : in     vl_logic_vector(31 downto 0);
        Stall           : in     vl_logic;
        WBDadoDeRetorno : in     vl_logic_vector(31 downto 0);
        WBEscreveReg    : in     vl_logic;
        WBMemParaReg    : in     vl_logic;
        Zero            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end PipelineInit_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Coproc_vlg_vec_tst is
end Coproc_vlg_vec_tst;

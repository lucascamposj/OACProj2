library verilog;
use verilog.vl_types.all;
entity IDEX_vlg_vec_tst is
end IDEX_vlg_vec_tst;

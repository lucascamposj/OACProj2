library verilog;
use verilog.vl_types.all;
entity Adder32_vlg_vec_tst is
end Adder32_vlg_vec_tst;

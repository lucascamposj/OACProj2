library verilog;
use verilog.vl_types.all;
entity controlPC_vlg_check_tst is
    port(
        JAL             : in     vl_logic;
        Jump            : in     vl_logic;
        JumpPC          : in     vl_logic_vector(31 downto 0);
        sampler_rx      : in     vl_logic
    );
end controlPC_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity mux1to2_vlg_check_tst is
    port(
        R               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux1to2_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Hazard_vlg_vec_tst is
end Hazard_vlg_vec_tst;

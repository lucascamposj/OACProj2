library verilog;
use verilog.vl_types.all;
entity controlALU_vlg_vec_tst is
end controlALU_vlg_vec_tst;

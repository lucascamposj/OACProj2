library IEEE;
use IEEE.STD_LOGIC_1164.all;
 
entity encoder32 is
 port(
 a : in STD_LOGIC_VECTOR(31 downto 0);
 b : out STD_LOGIC_VECTOR(5 downto 0)
 );
end encoder32;

architecture bhv of encoder32 is
begin
process(a)
begin
 case a is
  when "00000000000000000000000000000000" => b <= "000000"; 
  when "10000000000000000000000000000000" => b <= "000001"; 
  when "01000000000000000000000000000000" => b <= "000010"; 
  when "00100000000000000000000000000000" => b <= "000011"; 
  when "00010000000000000000000000000000" => b <= "000100"; 
  when "00001000000000000000000000000000" => b <= "000101"; 
  when "00000100000000000000000000000000" => b <= "000110"; 
  when "00000010000000000000000000000000" => b <= "000111"; 
  when "00000001000000000000000000000000" => b <= "001000"; 
  when "00000000100000000000000000000000" => b <= "001001"; 
  when "00000000010000000000000000000000" => b <= "001010"; 
  when "00000000001000000000000000000000" => b <= "001011"; 
  when "00000000000100000000000000000000" => b <= "001100"; 
  when "00000000000010000000000000000000" => b <= "001101"; 
  when "00000000000001000000000000000000" => b <= "001110"; 
  when "00000000000000100000000000000000" => b <= "001111"; 
  when "00000000000000010000000000000000" => b <= "010000"; 
  when "00000000000000001000000000000000" => b <= "010001"; 
  when "00000000000000000100000000000000" => b <= "010010"; 
  when "00000000000000000010000000000000" => b <= "010011"; 
  when "00000000000000000001000000000000" => b <= "010100"; 
  when "00000000000000000000100000000000" => b <= "010101"; 
  when "00000000000000000000010000000000" => b <= "010110"; 
  when "00000000000000000000001000000000" => b <= "010111"; 
  when "00000000000000000000000100000000" => b <= "011000"; 
  when "00000000000000000000000010000000" => b <= "011001"; 
  when "00000000000000000000000001000000" => b <= "011010"; 
  when "00000000000000000000000000100000" => b <= "011011"; 
  when "00000000000000000000000000010000" => b <= "011100"; 
  when "00000000000000000000000000001000" => b <= "011101"; 
  when "00000000000000000000000000000100" => b <= "011110"; 
  when "00000000000000000000000000000010" => b <= "011111"; 
  when "00000000000000000000000000000001" => b <= "100000";  
  when others => b <= "000000";
 end case;
end process;
end bhv;

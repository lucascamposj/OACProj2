library verilog;
use verilog.vl_types.all;
entity ula1bit_vlg_vec_tst is
end ula1bit_vlg_vec_tst;

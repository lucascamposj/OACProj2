library verilog;
use verilog.vl_types.all;
entity PipelineInit is
    port(
        OrigPC          : out    vl_logic;
        MEMZero         : out    vl_logic;
        clock           : in     vl_logic;
        DInstruction    : out    vl_logic_vector(31 downto 0);
        Flush           : out    vl_logic;
        Jump            : out    vl_logic;
        WBEscreveReg    : out    vl_logic;
        MEMReadValue    : out    vl_logic_vector(31 downto 0);
        MEMEscreveMem   : out    vl_logic;
        WBMemParaReg    : out    vl_logic;
        Stall           : out    vl_logic;
        clock2          : in     vl_logic;
        MEMnPC          : out    vl_logic_vector(31 downto 0);
        Zero            : out    vl_logic;
        ForwardA        : out    vl_logic_vector(1 downto 0);
        EXImm           : out    vl_logic_vector(5 downto 0);
        ForwardB        : out    vl_logic_vector(1 downto 0);
        EXopALU         : out    vl_logic_vector(2 downto 0);
        EXBranch        : out    vl_logic_vector(1 downto 0);
        outALU          : out    vl_logic_vector(31 downto 0);
        MEMBranch       : out    vl_logic_vector(1 downto 0);
        DJAL            : out    vl_logic;
        DJump           : out    vl_logic;
        DCtrlExtent     : out    vl_logic;
        DCtrlEscreveReg : out    vl_logic;
        DCtrlMemParaReg : out    vl_logic;
        DCtrlEscreveMem : out    vl_logic;
        DCtrlOrigALU    : out    vl_logic;
        ALUOperation    : out    vl_logic_vector(3 downto 0);
        BInstruction    : out    vl_logic_vector(31 downto 0);
        BPC             : out    vl_logic_vector(31 downto 0);
        BproxPC         : out    vl_logic_vector(31 downto 0);
        DCtrlBranch     : out    vl_logic_vector(1 downto 0);
        DCtrlcontrolJump: out    vl_logic_vector(1 downto 0);
        DCtrlopALU      : out    vl_logic_vector(2 downto 0);
        DCtrlRegDst     : out    vl_logic_vector(1 downto 0);
        DJumpPC         : out    vl_logic_vector(31 downto 0);
        DRSDados0       : out    vl_logic_vector(31 downto 0);
        DRTDados1       : out    vl_logic_vector(31 downto 0);
        EXHIGH          : out    vl_logic_vector(31 downto 0);
        EXLOW           : out    vl_logic_vector(31 downto 0);
        EXULAA          : out    vl_logic_vector(31 downto 0);
        EXULAB          : out    vl_logic_vector(31 downto 0);
        WBDadoDeRetorno : out    vl_logic_vector(31 downto 0)
    );
end PipelineInit;

library verilog;
use verilog.vl_types.all;
entity Equal_vlg_vec_tst is
end Equal_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity mux1to2_vlg_vec_tst is
end mux1to2_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity PipelineInit is
    port(
        OrigPC          : out    vl_logic;
        clock           : in     vl_logic;
        Flush           : out    vl_logic;
        Jump            : out    vl_logic;
        clock2          : in     vl_logic;
        MemReadValue    : out    vl_logic_vector(31 downto 0);
        MEMOutALU       : out    vl_logic_vector(31 downto 0);
        Stall           : out    vl_logic;
        notOpSignal     : out    vl_logic;
        JAL             : out    vl_logic;
        Zero            : out    vl_logic;
        ForwardA        : out    vl_logic_vector(1 downto 0);
        TreatedForwardB : out    vl_logic_vector(1 downto 0);
        ForwardB        : out    vl_logic_vector(1 downto 0);
        EXopALU         : out    vl_logic_vector(2 downto 0);
        EXBranch        : out    vl_logic_vector(1 downto 0);
        outALU          : out    vl_logic_vector(31 downto 0);
        MEMBranch       : out    vl_logic_vector(1 downto 0);
        WBMemPraReg     : out    vl_logic;
        ALUOperation    : out    vl_logic_vector(3 downto 0);
        atR             : out    vl_logic_vector(31 downto 0);
        BInstruction    : out    vl_logic_vector(31 downto 0);
        BPC             : out    vl_logic_vector(31 downto 0);
        EXULAA          : out    vl_logic_vector(31 downto 0);
        EXULAB          : out    vl_logic_vector(31 downto 0);
        RegA            : out    vl_logic_vector(31 downto 0);
        t0R             : out    vl_logic_vector(31 downto 0);
        t1R             : out    vl_logic_vector(31 downto 0);
        t2R             : out    vl_logic_vector(31 downto 0);
        t3R             : out    vl_logic_vector(31 downto 0);
        t4R             : out    vl_logic_vector(31 downto 0);
        t5R             : out    vl_logic_vector(31 downto 0);
        v0R             : out    vl_logic_vector(31 downto 0);
        WBDadoDeRetorno : out    vl_logic_vector(31 downto 0)
    );
end PipelineInit;

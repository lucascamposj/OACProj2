library verilog;
use verilog.vl_types.all;
entity mux1to2_vlg_sample_tst is
    port(
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        S               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end mux1to2_vlg_sample_tst;

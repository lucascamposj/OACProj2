library verilog;
use verilog.vl_types.all;
entity IFID_vlg_vec_tst is
end IFID_vlg_vec_tst;

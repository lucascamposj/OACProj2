library verilog;
use verilog.vl_types.all;
entity ShiftRight_vlg_vec_tst is
end ShiftRight_vlg_vec_tst;
